module top;
  initial begin
    $display("Hello PCIE UVM");
  end
endmodule
