interface pcie_tl_rc_intf(input bit clk,rst); 
logic[31:0] data;
    endinterface
