typedef uvm_sequencer#(pcie_tl_rc_mem_seq_item_pkg) pcie_tl_rc_sequencer;
